module decimal_to_bit (
        input [3:0] input,
        output pin 1,
        output pin 2,
        output pin 3,
        output pin 4,
        output pin 5,
        output pin 6,
        output pin 8
    );

    





endmodule